module my_module
  #(
    parameter integer MY_PARAM_0 = 0,
    parameter integer MY_PARAM_1 = 1,
    parameter integer MY_PARAM_2 = 2
    )
  (
   input wire clk,
   input wire rst,

   output reg A,
   output wire [7:0] B,
   output wire [(MY_PARAM_0-MY_PARAM_1)+MY_PARAM_2+1:0] C
   );

   //rest gets ignored for now!
   wire                        test;

endmodule
